

module Core (
    input wire clk,
    input wire startup
);






endmodule